module MUX_2to1();

endmodule